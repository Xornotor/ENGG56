module Semaforo (a, b, c, d, n_s, l_o);
input a, b, c, d;
output reg n_s, l_o;

endmodule