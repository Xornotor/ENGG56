module FSM ();

endmodule